/**************************************
@ filename    : print_pkg.sv
@ author      : yyrwkk
@ create time : 2025/06/15 23:02:25
@ version     : v1.0.0
**************************************/
package print_pkg;

function void show_pass();
begin: pass
    $display("pwd: %m");
    $display(".----------------.  .----------------.  .----------------.  .----------------. " ); 
    $display("| .--------------. || .--------------. || .--------------. || .--------------. |");
    $display("| |   ______     | || |      __      | || |    _______   | || |    _______   | |");
    $display("| |  |_   __ \\   | || |     /  \\     | || |   /  ___  |  | || |   /  ___  |  | |");
    $display("| |    | |__) |  | || |    / /\\ \\    | || |  |  (__ \\_|  | || |  |  (__ \\_|  | |");
    $display("| |    |  ___/   | || |   / ____ \\   | || |   '.___`-.   | || |   '.___`-.   | |");
    $display("| |   _| |_      | || | _/ /    \\ \\_ | || |  |`\\____) |  | || |  |`\\____) |  | |");
    $display("| |  |_____|     | || ||____|  |____|| || |  |_______.'  | || |  |_______.'  | |");
    $display("| |              | || |              | || |              | || |              | |");
    $display("| '--------------' || '--------------' || '--------------' || '--------------' |");
    $display("'----------------'  '----------------'  '----------------'  '----------------' " );   
    $display("time: %0t",$time );
end
endfunction

function void show_fail();
begin: fail
    $display("pwd: %m");
    $display(".----------------.  .----------------.  .----------------.  .----------------. " ); 
    $display("| .--------------. || .--------------. || .--------------. || .--------------. |");
    $display("| |  _________   | || |      __      | || |     _____    | || |   _____      | |");
    $display("| | |_   ___  |  | || |     /  \\     | || |    |_   _|   | || |  |_   _|     | |");
    $display("| |   |  _|      | || |   / ____ \\   | || |      | |     | || |    | |   _   | |");
    $display("| |  _| |_       | || | _/ /    \\ \\_ | || |     _| |_    | || |   _| |__/ |  | |");
    $display("| | |_____|      | || ||____|  |____|| || |    |_____|   | || |  |________|  | |");
    $display("| |              | || |              | || |              | || |              | |");
    $display("| '--------------' || '--------------' || '--------------' || '--------------' |");
    $display("'----------------'  '----------------'  '----------------'  '----------------' " );
    $display("time: %0t",$time );
end
endfunction

endpackage 